library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity NAND_GATE is
	Port
	(
		A : in STD_LOGIC; -- INPUT A
		B : in STD_LOGIC; -- INPUT B
		Y : out STD_LOGIC -- OUTPUT Y
	);
end NAND_GATE;
architecture Behavior of NAND_GATE is begin
	Y <= A NAND B;
end Behavior;
